//: version "1.8.3"

module OR(X, B, A);
//: interface  /sz:(40, 40) /bd:[ Li0>A(10/40) Li1>B(26/40) Ro0<X(20/40) ]
input B;    //: /sn:0 /dp:1 {0}(277,310)(220,310){1}
//: {2}(218,308)(218,101)(333,101){3}
//: {4}(216,310)(179,310)(179,269)(171,269){5}
output X;    //: /sn:0 {0}(347,110)(347,210){1}
//: {2}(349,212)(365,212){3}
//: {4}(369,212)(496,212){5}
//: {6}(367,214)(367,302){7}
//: {8}(345,212)(291,212)(291,302){9}
input A;    //: /sn:0 /dp:1 {0}(353,310)(333,310)(333,188)(206,188){1}
//: {2}(204,186)(204,52)(333,52){3}
//: {4}(202,188)(170,188){5}
supply0 w0;    //: /sn:0 {0}(309,28)(309,18)(347,18)(347,44){1}
supply1 w2;    //: /sn:0 {0}(367,319)(367,371)(324,371){1}
//: {2}(322,369)(322,353){3}
//: {4}(320,371)(291,371)(291,319){5}
wire w7;    //: /sn:0 /dp:1 {0}(347,61)(347,93){1}
//: enddecls

  nmos g4 (.Z(w2), .S0(X), .G0(A));   //: @(361,310) /sn:0 /w:[ 0 7 0 ]
  //: joint g8 (w2) @(322, 371) /w:[ 1 2 4 -1 ]
  nmos g3 (.Z(w2), .S0(X), .G0(B));   //: @(285,310) /sn:0 /w:[ 5 9 0 ]
  //: joint g13 (X) @(347, 212) /w:[ 2 1 8 -1 ]
  //: output g2 (X) @(493,212) /sn:0 /w:[ 5 ]
  //: input g1 (B) @(169,269) /sn:0 /w:[ 5 ]
  //: supply0 g11 (w0) @(309,34) /sn:0 /w:[ 0 ]
  //: joint g10 (B) @(218, 310) /w:[ 1 2 4 -1 ]
  pmos g6 (.Z(w7), .S0(X), .G0(B));   //: @(341,101) /sn:0 /w:[ 1 0 3 ]
  //: supply1 g7 (w2) @(333,353) /sn:0 /w:[ 3 ]
  //: joint g9 (A) @(204, 188) /w:[ 1 2 4 -1 ]
  pmos g5 (.Z(w0), .S0(w7), .G0(A));   //: @(341,52) /sn:0 /w:[ 1 0 3 ]
  //: comment g14 /dolink:0 /link:"" @(467,76) /sn:0
  //: /line:"OR gate: 4 transistors"
  //: /end
  //: input g0 (A) @(168,188) /sn:0 /w:[ 5 ]
  //: joint g12 (X) @(367, 212) /w:[ 4 -1 3 6 ]

endmodule

module XOR(X, B, A);
//: interface  /sz:(40, 40) /bd:[ Li0>A(9/40) Li1>B(26/40) Ro0<X(17/40) ]
input B;    //: /sn:0 {0}(167,242)(254,242){1}
//: {2}(258,242)(266,242){3}
//: {4}(256,240)(256,197)(265,197){5}
output X;    //: /sn:0 {0}(461,202)(520,202){1}
input A;    //: /sn:0 /dp:1 {0}(265,182)(245,182){1}
//: {2}(241,182)(169,182){3}
//: {4}(243,184)(243,225)(266,225){5}
wire w0;    //: /sn:0 {0}(333,236)(308,236){1}
wire w1;    //: /sn:0 {0}(375,237)(409,237)(409,208)(419,208){1}
wire w2;    //: /sn:0 {0}(307,191)(419,191){1}
//: enddecls

  AND g4 (.A(A), .B(B), .X(w0));   //: @(267, 217) /sz:(40, 40) /sn:0 /p:[ Li0>5 Li1>3 Ro0<1 ]
  AND g8 (.A(w2), .B(w1), .X(X));   //: @(420, 183) /sz:(40, 40) /sn:0 /p:[ Li0>1 Li1>1 Ro0<0 ]
  OR g3 (.A(A), .B(B), .X(w2));   //: @(266, 171) /sz:(40, 40) /sn:0 /p:[ Li0>0 Li1>5 Ro0<0 ]
  //: output g2 (X) @(517,202) /sn:0 /w:[ 1 ]
  //: input g1 (B) @(165,242) /sn:0 /w:[ 0 ]
  //: joint g6 (B) @(256, 242) /w:[ 2 4 1 -1 ]
  NOT g7 (.A(w0), .X(w1));   //: @(334, 219) /sz:(40, 40) /sn:0 /p:[ Li0>0 Ro0<0 ]
  //: comment g9 /dolink:0 /link:"" @(421,89) /sn:0
  //: /line:"XOR gate: 14 transistors"
  //: /end
  //: joint g5 (A) @(243, 182) /w:[ 1 -1 2 4 ]
  //: input g0 (A) @(167,182) /sn:0 /w:[ 3 ]

endmodule

module ADD8(R, X, C, B, A);
//: interface  /sz:(40, 40) /bd:[ Ti0>C(19/40) Li0>A[7:0](10/40) Li1>B[7:0](30/40) Bo0<R(20/40) Ro0<X[7:0](22/40) ]
input [7:0] B;    //: /sn:0 {0}(-18,594)(49,594){1}
//: {2}(50,594)(68,594){3}
//: {4}(69,594)(90,594){5}
//: {6}(91,594)(109,594){7}
//: {8}(110,594)(131,594){9}
//: {10}(132,594)(154,594){11}
//: {12}(155,594)(177,594){13}
//: {14}(178,594)(194,594){15}
//: {16}(195,594)(222,594){17}
output [7:0] X;    //: /sn:0 {0}(652,276)(536,276){1}
input [7:0] A;    //: /sn:0 {0}(-9,56)(77,56){1}
//: {2}(78,56)(100,56){3}
//: {4}(101,56)(120,56){5}
//: {6}(121,56)(142,56){7}
//: {8}(143,56)(166,56){9}
//: {10}(167,56)(186,56){11}
//: {12}(187,56)(203,56){13}
//: {14}(204,56)(219,56){15}
//: {16}(220,56)(247,56){17}
output R;    //: /sn:0 {0}(351,565)(351,595)(411,595){1}
input C;    //: /sn:0 {0}(317,34)(361,34)(361,72){1}
wire w6;    //: /sn:0 {0}(178,589)(178,162)(339,162){1}
wire w32;    //: /sn:0 {0}(101,60)(101,466)(332,466){1}
wire w7;    //: /sn:0 {0}(204,60)(204,146)(339,146){1}
wire w16;    //: /sn:0 {0}(132,589)(132,289)(336,289){1}
wire w15;    //: /sn:0 {0}(358,264)(358,243){1}
wire w38;    //: /sn:0 {0}(530,241)(435,241)(435,541)(373,541){1}
wire w0;    //: /sn:0 {0}(530,311)(483,311)(483,90)(382,90){1}
wire w3;    //: /sn:0 {0}(530,301)(475,301)(475,155)(381,155){1}
wire w37;    //: /sn:0 {0}(78,60)(78,532)(331,532){1}
wire w21;    //: /sn:0 {0}(110,589)(110,353)(334,353){1}
wire w31;    //: /sn:0 {0}(69,589)(69,482)(332,482){1}
wire w28;    //: /sn:0 {0}(530,261)(453,261)(453,411)(375,411){1}
wire w20;    //: /sn:0 {0}(356,328)(356,306){1}
wire w36;    //: /sn:0 {0}(50,589)(50,548)(331,548){1}
wire w23;    //: /sn:0 {0}(530,271)(459,271)(459,346)(376,346){1}
wire w1;    //: /sn:0 {0}(195,589)(195,97)(340,97){1}
wire w25;    //: /sn:0 {0}(354,393)(354,370){1}
wire w35;    //: /sn:0 {0}(352,523)(352,499){1}
wire w18;    //: /sn:0 {0}(530,281)(387,281)(387,282)(378,282){1}
wire w30;    //: /sn:0 {0}(353,457)(353,435){1}
wire w17;    //: /sn:0 {0}(167,60)(167,273)(336,273){1}
wire w22;    //: /sn:0 {0}(143,60)(143,337)(334,337){1}
wire w2;    //: /sn:0 {0}(220,60)(220,81)(340,81){1}
wire w11;    //: /sn:0 {0}(155,589)(155,226)(338,226){1}
wire w12;    //: /sn:0 {0}(187,60)(187,210)(338,210){1}
wire w10;    //: /sn:0 {0}(359,201)(359,179){1}
wire w27;    //: /sn:0 {0}(121,60)(121,402)(333,402){1}
wire w13;    //: /sn:0 {0}(530,291)(467,291)(467,221)(380,221){1}
wire w5;    //: /sn:0 {0}(360,137)(360,114){1}
wire w33;    //: /sn:0 {0}(530,251)(444,251)(444,475)(374,475){1}
wire w26;    //: /sn:0 {0}(91,589)(91,418)(333,418){1}
//: enddecls

  //: output g4 (R) @(408,595) /sn:0 /w:[ 1 ]
  BADD g8 (.C(w15), .A(w17), .B(w16), .R(w20), .X(w18));   //: @(337, 265) /sz:(40, 40) /sn:0 /p:[ Ti0>0 Li0>1 Li1>1 Bo0<1 Ro0<1 ]
  //: output g3 (X) @(649,276) /sn:0 /w:[ 0 ]
  tran g13(.Z(w2), .I(A[0]));   //: @(220,54) /sn:0 /R:1 /w:[ 0 15 16 ] /ss:1
  //: input g2 (C) @(315,34) /sn:0 /w:[ 0 ]
  //: input g1 (B) @(-20,594) /sn:0 /w:[ 0 ]
  BADD g11 (.C(w30), .A(w32), .B(w31), .R(w35), .X(w33));   //: @(333, 458) /sz:(40, 40) /sn:0 /p:[ Ti0>0 Li0>1 Li1>1 Bo0<1 Ro0<1 ]
  tran g16(.Z(w17), .I(A[3]));   //: @(167,54) /sn:0 /R:1 /w:[ 0 9 10 ] /ss:1
  BADD g10 (.C(w25), .A(w27), .B(w26), .R(w30), .X(w28));   //: @(334, 394) /sz:(40, 40) /sn:0 /p:[ Ti0>0 Li0>1 Li1>1 Bo0<1 Ro0<1 ]
  tran g28(.Z(w36), .I(B[7]));   //: @(50,592) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:0
  tran g19(.Z(w32), .I(A[6]));   //: @(101,54) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  tran g27(.Z(w31), .I(B[6]));   //: @(69,592) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:0
  BADD g6 (.C(w5), .A(w7), .B(w6), .R(w10), .X(w3));   //: @(340, 138) /sz:(40, 40) /sn:0 /p:[ Ti0>0 Li0>1 Li1>1 Bo0<1 Ro0<1 ]
  BADD g7 (.C(w10), .A(w12), .B(w11), .R(w15), .X(w13));   //: @(339, 202) /sz:(40, 40) /sn:0 /p:[ Ti0>0 Li0>1 Li1>1 Bo0<1 Ro0<1 ]
  BADD g9 (.C(w20), .A(w22), .B(w21), .R(w25), .X(w23));   //: @(335, 329) /sz:(40, 40) /sn:0 /p:[ Ti0>0 Li0>1 Li1>1 Bo0<1 Ro0<1 ]
  tran g15(.Z(w12), .I(A[2]));   //: @(187,54) /sn:0 /R:1 /w:[ 0 11 12 ] /ss:1
  tran g20(.Z(w37), .I(A[7]));   //: @(78,54) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  tran g17(.Z(w22), .I(A[4]));   //: @(143,54) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1
  tran g25(.Z(w21), .I(B[4]));   //: @(110,592) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:0
  concat g29 (.I0(w0), .I1(w3), .I2(w13), .I3(w18), .I4(w23), .I5(w28), .I6(w33), .I7(w38), .Z(X));   //: @(535,276) /sn:0 /w:[ 0 0 0 0 0 0 0 0 1 ] /dr:0
  BADD g5 (.C(C), .A(w2), .B(w1), .R(w5), .X(w0));   //: @(341, 73) /sz:(40, 40) /sn:0 /p:[ Ti0>1 Li0>1 Li1>1 Bo0<1 Ro0<1 ]
  tran g14(.Z(w7), .I(A[1]));   //: @(204,54) /sn:0 /R:1 /w:[ 0 13 14 ] /ss:1
  tran g21(.Z(w1), .I(B[0]));   //: @(195,592) /sn:0 /R:1 /w:[ 0 15 16 ] /ss:0
  tran g24(.Z(w16), .I(B[3]));   //: @(132,592) /sn:0 /R:1 /w:[ 0 9 10 ] /ss:0
  tran g23(.Z(w11), .I(B[2]));   //: @(155,592) /sn:0 /R:1 /w:[ 0 11 12 ] /ss:0
  //: input g0 (A) @(-11,56) /sn:0 /w:[ 0 ]
  tran g22(.Z(w6), .I(B[1]));   //: @(178,592) /sn:0 /R:1 /w:[ 0 13 14 ] /ss:0
  tran g26(.Z(w26), .I(B[5]));   //: @(91,592) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:0
  BADD g12 (.C(w35), .A(w37), .B(w36), .R(R), .X(w38));   //: @(332, 524) /sz:(40, 40) /sn:0 /p:[ Ti0>0 Li0>1 Li1>1 Bo0<0 Ro0<1 ]
  tran g18(.Z(w27), .I(A[5]));   //: @(121,54) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1
  //: comment g30 /dolink:0 /link:"" @(536,73) /sn:0
  //: /line:"ADD8 gate: 320 transistors"
  //: /end

endmodule

module BADD(R, X, C, B, A);
//: interface  /sz:(40, 40) /bd:[ Ti0>C(20/40) Li0>A(8/40) Li1>B(24/40) Bo0<R(19/40) Ro0<X(17/40) ]
input B;    //: /sn:0 {0}(174,203)(196,203){1}
//: {2}(200,203)(226,203)(226,172)(230,172){3}
//: {4}(198,205)(198,332)(261,332){5}
output X;    //: /sn:0 {0}(339,206)(566,206)(566,180)(577,180){1}
input A;    //: /sn:0 {0}(174,155)(211,155){1}
//: {2}(215,155)(230,155){3}
//: {4}(213,157)(213,317)(261,317){5}
output R;    //: /sn:0 {0}(578,224)(568,224)(568,295)(410,295){1}
input C;    //: /sn:0 /dp:1 {0}(172,244)(236,244)(236,213)(274,213){1}
//: {2}(278,213)(297,213){3}
//: {4}(276,215)(276,279)(300,279){5}
wire w6;    //: /sn:0 {0}(303,328)(358,328)(358,301)(368,301){1}
wire w3;    //: /sn:0 {0}(342,270)(358,270)(358,287)(368,287){1}
wire w1;    //: /sn:0 {0}(297,198)(285,198){1}
//: {2}(283,196)(283,163)(272,163){3}
//: {4}(283,200)(283,262)(300,262){5}
//: enddecls

  //: output g4 (R) @(575,224) /sn:0 /w:[ 0 ]
  AND g8 (.A(A), .B(B), .X(w6));   //: @(262, 309) /sz:(40, 40) /sn:0 /p:[ Li0>5 Li1>5 Ro0<0 ]
  //: output g3 (X) @(574,180) /sn:0 /w:[ 1 ]
  //: joint g13 (C) @(276, 213) /w:[ 2 -1 1 4 ]
  //: input g2 (C) @(170,244) /sn:0 /w:[ 0 ]
  //: input g1 (B) @(172,203) /sn:0 /w:[ 0 ]
  //: joint g11 (B) @(198, 203) /w:[ 2 -1 1 4 ]
  //: joint g10 (A) @(213, 155) /w:[ 2 -1 1 4 ]
  XOR g6 (.A(w1), .B(C), .X(X));   //: @(298, 189) /sz:(40, 40) /sn:0 /p:[ Li0>0 Li1>3 Ro0<0 ]
  AND g7 (.A(w1), .B(C), .X(w3));   //: @(301, 254) /sz:(40, 40) /sn:0 /p:[ Li0>5 Li1>5 Ro0<0 ]
  OR g9 (.A(w3), .B(w6), .X(R));   //: @(369, 275) /sz:(40, 40) /sn:0 /p:[ Li0>1 Li1>1 Ro0<1 ]
  XOR g5 (.A(A), .B(B), .X(w1));   //: @(231, 146) /sz:(40, 40) /sn:0 /p:[ Li0>3 Li1>3 Ro0<3 ]
  //: comment g14 /dolink:0 /link:"" @(474,55) /sn:0
  //: /line:"BADD Gate: 40 transistors."
  //: /end
  //: input g0 (A) @(172,155) /sn:0 /w:[ 0 ]
  //: joint g12 (w1) @(283, 198) /w:[ 1 2 -1 4 ]

endmodule

module main;    //: root_module
wire [7:0] w4;    //: /sn:0 {0}(399,149)(399,215)(332,215){1}
wire w0;    //: /sn:0 {0}(388,256)(388,266)(311,266)(311,234){1}
wire w1;    //: /sn:0 {0}(292,115)(310,115)(310,192){1}
wire [7:0] w2;    //: /sn:0 {0}(186,172)(186,219)(290,219){1}
wire [7:0] w5;    //: /sn:0 {0}(102,172)(102,203)(290,203){1}
//: enddecls

  led g4 (.I(w0));   //: @(388,249) /sn:0 /w:[ 0 ] /type:0
  //: switch g3 (w1) @(275,115) /sn:0 /w:[ 0 ] /st:0
  //: dip g2 (w2) @(186,162) /sn:0 /w:[ 0 ] /st:63
  //: dip g1 (w5) @(102,162) /sn:0 /w:[ 0 ] /st:208
  led g5 (.I(w4));   //: @(399,142) /sn:0 /w:[ 0 ] /type:2
  ADD8 g0 (.C(w1), .A(w5), .B(w2), .R(w0), .X(w4));   //: @(291, 193) /sz:(40, 40) /sn:0 /p:[ Ti0>1 Li0>1 Li1>1 Bo0<1 Ro0<1 ]

endmodule

module NOT(X, A);
//: interface  /sz:(40, 40) /bd:[ Li0>A(17/40) Ro0<X(18/40) ]
supply1 w6;    //: /sn:0 {0}(339,135)(339,159){1}
output X;    //: /sn:0 /dp:1 {0}(339,229)(339,203){1}
//: {2}(341,201)(377,201){3}
//: {4}(339,199)(339,176){5}
supply0 w7;    //: /sn:0 {0}(339,271)(339,246){1}
input A;    //: /sn:0 /dp:1 {0}(325,167)(269,167)(269,203){1}
//: {2}(267,205)(150,205){3}
//: {4}(269,207)(269,237)(325,237){5}
//: enddecls

  //: supply1 g4 (w6) @(350,135) /sn:0 /w:[ 0 ]
  //: comment g8 /dolink:0 /link:"" @(424,77) /sn:0
  //: /line:"Not Gate: 2 transistors"
  //: /end
  pmos g3 (.Z(w6), .S0(X), .G0(A));   //: @(333,167) /sn:0 /w:[ 1 5 0 ]
  nmos g2 (.Z(w7), .S0(X), .G0(A));   //: @(333,237) /sn:0 /w:[ 1 0 5 ]
  //: output g1 (X) @(374,201) /sn:0 /w:[ 3 ]
  //: joint g6 (A) @(269, 205) /w:[ -1 1 2 4 ]
  //: joint g7 (X) @(339, 201) /w:[ 2 4 -1 1 ]
  //: supply0 g5 (w7) @(339,277) /sn:0 /w:[ 0 ]
  //: input g0 (A) @(148,205) /sn:0 /w:[ 3 ]

endmodule

module AND(X, B, A);
//: interface  /sz:(40, 40) /bd:[ Li0>A(8/40) Li1>B(25/40) Ro0<X(19/40) ]
input B;    //: /sn:0 {0}(181,280)(227,280){1}
//: {2}(231,280)(327,280)(327,159)(343,159){3}
//: {4}(229,282)(229,383)(302,383){5}
output X;    //: /sn:0 {0}(316,323)(316,265){1}
//: {2}(318,263)(355,263){3}
//: {4}(359,263)(505,263){5}
//: {6}(357,261)(357,168){7}
//: {8}(314,263)(306,263)(306,169){9}
input A;    //: /sn:0 {0}(177,218)(253,218){1}
//: {2}(255,216)(255,160)(292,160){3}
//: {4}(255,220)(255,331)(302,331){5}
supply0 w0;    //: /sn:0 {0}(306,152)(306,129)(355,129){1}
//: {2}(359,129)(401,129)(401,139){3}
//: {4}(357,131)(357,151){5}
supply1 w12;    //: /sn:0 {0}(262,404)(262,429)(316,429)(316,392){1}
wire w4;    //: /sn:0 {0}(316,375)(316,340){1}
//: enddecls

  nmos g4 (.Z(w12), .S0(w4), .G0(B));   //: @(310,383) /sn:0 /w:[ 1 0 5 ]
  //: joint g8 (A) @(255, 218) /w:[ -1 2 1 4 ]
  nmos g3 (.Z(w4), .S0(X), .G0(A));   //: @(310,331) /sn:0 /w:[ 1 0 5 ]
  //: joint g13 (X) @(316, 263) /w:[ 2 -1 8 1 ]
  //: output g2 (X) @(502,263) /sn:0 /w:[ 5 ]
  //: input g1 (B) @(179,280) /sn:0 /w:[ 0 ]
  //: joint g11 (w0) @(357, 129) /w:[ 2 -1 1 4 ]
  //: supply0 g10 (w0) @(401,145) /sn:0 /w:[ 3 ]
  pmos g6 (.Z(w0), .S0(X), .G0(B));   //: @(351,159) /sn:0 /w:[ 5 7 3 ]
  //: supply1 g7 (w12) @(273,404) /sn:0 /w:[ 0 ]
  //: joint g9 (B) @(229, 280) /w:[ 2 -1 1 4 ]
  pmos g5 (.Z(w0), .S0(X), .G0(A));   //: @(300,160) /sn:0 /w:[ 0 9 3 ]
  //: comment g14 /dolink:0 /link:"" @(471,72) /sn:0
  //: /line:"AND gate: 4 transistors"
  //: /end
  //: input g0 (A) @(175,218) /sn:0 /w:[ 0 ]
  //: joint g12 (X) @(357, 263) /w:[ 4 6 3 -1 ]

endmodule
